module ram_char (
	input  [6:0]   raddr,
	output [511:0] rdata
);

reg [511:0] ram[23:0];
assign rdata = ram[raddr];

initial
begin
	ram[0] = 512'h00000000000000000000000003C006200C30181818181808300C300C300C300C300C300C300C300C300C300C1808181818180C30062003C00000000000000000;
	ram[1] = 512'h000000000000000000000000008001801F800180018001800180018001800180018001800180018001800180018001800180018003C01FF80000000000000000;
	ram[2] = 512'h00000000000000000000000007E008381018200C200C300C300C000C001800180030006000C0018003000200040408041004200C3FF83FF80000000000000000;
	ram[3] = 512'h00000000000000000000000007C018603030301830183018001800180030006003C0007000180008000C000C300C300C30083018183007C00000000000000000;
	ram[4] = 512'h0000000000000000000000000060006000E000E0016001600260046004600860086010603060206040607FFC0060006000600060006003FC0000000000000000;
	ram[5] = 512'h0000000000000000000000000FFC0FFC10001000100010001000100013E0143018181008000C000C000C000C300C300C20182018183007C00000000000000000;
	ram[6] = 512'h00000000000000000000000001E006180C180818180010001000300033E0363038183808300C300C300C300C300C180C18080C180E3003E00000000000000000;
	ram[7] = 512'h0000000000000000000000001FFC1FFC100830102010202000200040004000400080008001000100010001000300030003000300030003000000000000000000;
	ram[8] = 512'h00000000000000000000000007E00C301818300C300C300C380C38081E180F2007C018F030783038601C600C600C600C600C3018183007C00000000000000000;
	ram[9] = 512'h00000000000000000000000007C01820301030186008600C600C600C600C600C701C302C186C0F8C000C0018001800103030306030C00F800000000000000000;

	ram[10] = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
	
	ram[11] = 512'h00000000000000000000000000000000000000000000000000000000000000007FFE000000000000000000000000000000000000000000000000000000000000;
	ram[12] = 512'h00000000000000000000000020001000080004000200010000800040002000100008000800100020004000800100020004000800100020000000000000000000;
	ram[13] = 512'h00000000000000000000000000000000000000000000000000003E7C0C100E100620034003400180018001C0026004600430081818187C7E0000000000000000;

	ram[14] = 512'h000000000000000000000000000000000000000000000000000007E01830301830183018003807D81C183018601860186018601930791F8E0000000000000000;
	ram[15] = 512'h000000000000000000000800780018001800180018001800180019E01A381C181C0C180C180C180C180C180C180C180C18081C181C3013E00000000000000000;
	ram[16] = 512'h000000000000000000000000000000000000000000000000000003C00C3008181808300C300C300C3FFC300030003000180418080E1803E00000000000000000;
	ram[17] = 512'h000000000000000000000000000000000000000000000000000003EE0C36081818181818181808180C300FE0180018001FC00FF8181C300C300C300C181807E0;
	ram[18] = 512'h000000000000000000000800780018001800180018001800180019E01A301C18181818181818181818181818181818181818181818187E7E0000000000000000;
	ram[19] = 512'h000000000000000000000000018003C0018000000000000000801F8001800180018001800180018001800180018001800180018001801FF80000000000000000;
	ram[20] = 512'h0000000000000000000000801F80018001800180018001800180018001800180018001800180018001800180018001800180018001801FF80000000000000000;
	ram[21] = 512'h000000000000000000000000000000000000000000000000000009E07A301C18181818181818181818181818181818181818181818187E7E0000000000000000;
	ram[22] = 512'h000000000000000000000000000000000000000000000000000003C00C3008181818100C300C300C300C300C300C300C181818180C3003C00000000000000000;
	ram[23] = 512'h0000000000000000000000000000000000000000000000000000061C7E660686078007000600060006000600060006000600060006007FE00000000000000000;
end

endmodule






/////////////////// DdrRdCtrl ///////////////////////////////////
/**********************************************************
  Function Description:

  Establishment : Richard Zhu
  Create date   : 2020-01-09
  Versions      : V0.1
  Revision of records:
  Ver0.1

**********************************************************/
module  DdrRdCtrl #(
  parameter   TCo_C           = 1,

  parameter   AXI_RD_ID       = 8'ha5             ,
  parameter  	AXI_ID_WIDTH		= 8									,
  parameter   AXI_DATA_WIDTH  = 256               ,

  localparam  AXI_BYTE_NUMBER = AXI_DATA_WIDTH/8  ,
  localparam  AXI_DATA_SIZE   = $clog2(AXI_BYTE_NUMBER) ,  
  
  localparam  ADW_C           = AXI_DATA_WIDTH    ,
  localparam  ABN_C           = AXI_BYTE_NUMBER   


)
(
  /////////////////////////////////////////////////////////

  //Define Port
  /////////////////////////////////////////////////////////
  //System Signal
  input   wire		      	SysClk    ,     //System Clock
  input   wire		      	Reset_N   ,     //System Reset

  /////////////////////////////////////////////////////////
  //Operate Control & State
  input               		RamRdStart  , //(I)[DdrRdCtrl]Ram Read Start
  output  reg       		RamRdEnd    , //(O)[DdrRdCtrl]Ram Read End
  output  reg [     31:0] 	RamRdAddr   , //(O)[DdrRdCtrl]Ram Read Addrdss
  output  reg        		RamRdDAva   , //(O)[DdrRdCtrl]Ram Read Available
  output  reg           	RamRdBusy   , //(O)Ram Read Busy
  output              		RamRdALoad  , //(O)Ram Read Address Load
  output  reg [ADW_C-1:0] 	RamRdData   , //(O)[DdrRdCtrl]Ram Read Data

  /////////////////////////////////////////////////////////
  //Config DDR & AXI Operate Parameter
  input   [     31:0] 		CfgRdAddr   , //(I)[DdrRdCtrl]Config Read Start Address
  input   [      7:0] 		CfgRdBLen   , //(I)[DdrRdCtrl]Config Read Burst Length

  /////////////////////////////////////////////////////////
  //Axi4 Read Address & Data Bus
  output  [AXI_ID_WIDTH-1:0] 		ARID        , //(I)[RdAddr]Read address ID. This signal is the identification tag for the read address group of signals.
  output  [     31:0] 		ARADDR      , //(I)[RdAddr]Read address. The read address gives the address of the first transfer in a read burst transaction.
  output  [      7:0] 		ARLEN       , //(I)[RdAddr]Burst length. This signal indicates the exact number of transfers in a burst.
  output  [      2:0] 		ARSIZE      , //(I)[RdAddr]Burst size. This signal indicates the size of each transfer in the burst.
  output  [      1:0] 		ARBURST     , //(I)[RdAddr]Burst type. The burst type and the size information determine how the address for each transfer within the burst is calculated.
  output  [      1:0] 		ARLOCK      , //(I)[RdAddr]Lock type. This signal provides additional information about the atomic characteristics of the transfer.
  output              		ARVALID     , //(I)[RdAddr]Read address valid. This signal indicates that the channel is signaling valid read address and control information.
  input               		ARREADY     , //(O)[RdAddr]Read address ready. This signal indicates that the slave is ready to accept an address and associated control signals.
  /////////////       		       
  input   [AXI_ID_WIDTH-1:0] 		RID         , //(O)[RdData]Read ID tag. This signal is the identification tag for the read data group of signals generated by the slave.
  input   [      1:0] 		RRESP       , //(O)[RdData]Read response. This signal indicates the status of the read transfer.
  input               		RLAST       , //(O)[RdData]Read last. This signal indicates the last transfer in a read burst.
  input               		RVALID      , //(O)[RdData]Read valid. This signal indicates that the channel is signaling the required read data.
  output              		RREADY      , //(I)[RdData]Read ready. This signal indicates that the master can accept the read data and response information.
  input   [ADW_C-1:0] 		RDATA        //(O)[RdData]Read data.

);

  //Define  Parameter
  /////////////////////////////////////////////////////////
  reg   [7 :0]  RdBurstLen  = 8'h0;
  reg   [31:0]  RdStartAddr = 32'h0;
  reg     		AddrValid = 1'h0; //(I)[RdAddr]Read address valid. This signal indicates that the channel is signaling valid read address and control information.
  reg 	  	  	DataRdEndReg;
  reg 	[7:0] 	RdBurstCnt      = 8'h0;
  reg 	      	DataRdLastFlag  = 1'h0;
  reg 	[7:0] 	DataRdTimeOut   = 8'hff ;
  reg 	      	DataRdReadyClr  = 1'h0  ;
  reg   		DataRdAddrAva     = 1'h0;
  reg   		DataRdNextBrst    = 1'h0;
  reg   		DataRdStart       = 1'h0;
  reg   		DataRdReady = 1'h0; 

  /////////////////////////////////////////////////////////
  /////////////////////////////////////////////////////////
  assign  ARID    = AXI_RD_ID     ; //(I)[RdAddr]Read address ID. This signal is the identification tag for the read address group of signals.
  assign  ARADDR  = RdStartAddr   ; //(I)[RdAddr]Read address. The read address gives the address of the first transfer in a read burst transaction.
  assign  ARLEN   = RdBurstLen    ; //(I)[RdAddr]Burst length. This signal indicates the exact number of transfers in a burst.
  assign  ARSIZE  = AXI_DATA_SIZE ; //(I)[RdAddr]Burst size. This signal indicates the size of each transfer in the burst.
  assign  ARBURST = 2'b01         ; //(I)[RdAddr]Burst type. The burst type and the size information determine how the address for each transfer within the burst is calculated.
  assign  ARLOCK  = 2'h00         ; //(I)[RdAddr]Lock type. This signal provides additional information about the atomic characteristics of the transfer.
  assign  ARVALID = AddrValid     ; //(I)[RdAddr]Read address valid. This signal indicates that the channel is signaling valid read address and control information.
//  assign  RID 		= AXI_RD_ID     ; //(O)[RdData]Read ID tag. This signal is the identification tag for the read data group of signals generated by the slave.
  wire  [     1:0]   DataRdResp  = RRESP   ; //(O)[RdData]Read response. This signal indicates the status of the read transfer.
  wire               DataRdLast  = RLAST   ; //(O)[RdData]Read last. This signal indicates the last transfer in a read burst.
  wire               DataRdValid = RVALID  ; //(O)[RdData]Read valid. This signal indicates that the channel is signaling the required read data.
  wire  [ADW_C-1:0]  DataRdData  = RDATA   ; //(O)[RdData]Read data.
  assign  RREADY  = DataRdReady ; //(I)[RdData]Read ready. This signal indicates that the master can accept the read data and response information.

//1111111111111111111111111111111111111111111111111111111
//  Process AXI Operate Parameter
//  Input��
//  output��
//***************************************************/

  /////////////////////////////////////////////////////////
  wire  AddrReady = ARREADY;

  /////////////////////////////////////////////////////////
  

  always @( posedge SysClk)   if(RamRdStart)  RdBurstLen    <=   CfgRdBLen;
  always @( posedge SysClk)   if(RamRdStart)  RdStartAddr   <=   CfgRdAddr;

  /////////////////////////////////////////////////////////
  
  always @( posedge SysClk or negedge Reset_N)
  begin
    if (!Reset_N)         AddrValid <=  1'h0;
    else if (RamRdStart)  AddrValid <=  1'h1;
    else if (AddrReady)   AddrValid <=  1'h0;
  end

  wire AddrRdEn = (AddrValid & AddrReady);

  
//1111111111111111111111111111111111111111111111111111111



//22222222222222222222222222222222222222222222222222222
  /////////////////////////////////////////////////////////
  

  wire  DataRdEn    = DataRdReady & DataRdValid;
  wire  DataRdEnd   = DataRdReady & DataRdValid & DataRdLast;

  /////////////////////////////////////////////////////////
  
  always @( posedge SysClk or negedge Reset_N)
  begin
    if (~Reset_N)       DataRdAddrAva <=  1'h0;
    else if (DataRdEnd) DataRdAddrAva <=  1'h0;
    else if (AddrRdEn)  DataRdAddrAva <=  DataRdReady;
  end

  always @( posedge SysClk)  DataRdNextBrst <=  (AddrRdEn | DataRdAddrAva ) & DataRdEnd;
  always @( posedge SysClk)  DataRdStart    <=  (AddrRdEn & (~DataRdReady)) | DataRdNextBrst;

  assign  RamRdALoad =  DataRdStart; //(O)Ram Read Address Load;

  /////////////////////////////////////////////////////////
  

  always @( posedge SysClk)
  begin
    if (DataRdValid)  DataRdTimeOut <=  8'hff;
    else              DataRdTimeOut <=  DataRdTimeOut - {7'h0, (|DataRdTimeOut)};
  end

  always @( posedge SysClk)  DataRdReadyClr <=  (DataRdTimeOut == 5'h1);

  /////////////////////////////////////////////////////////
  

  always @( posedge SysClk or negedge Reset_N)
  begin
    if (! Reset_N)          RdBurstCnt <=  8'h0;
    else if (DataRdStart)   RdBurstCnt <=  RdBurstLen;
    else if (DataRdEn)      RdBurstCnt <=  RdBurstCnt - {7'h0,(|RdBurstCnt)};
  end

  always @( posedge SysClk)
  begin
    if (DataRdStart)    DataRdLastFlag <=  (RdBurstLen == 8'h0);
    else if (DataRdEn)  DataRdLastFlag <=  (RdBurstCnt == 8'h1);
    else if (DataRdEnd) DataRdLastFlag <=  (RdBurstCnt == 8'h0);
  end

  wire  DataRdEndFlag = DataRdLastFlag & DataRdEn;

  /////////////////////////////////////////////////////////
  
  
  always @( posedge SysClk)  DataRdEndReg <=  DataRdEnd;
  
  
  /////////////////////////////////////////////////////////
  always @( posedge SysClk )//or negedge Reset_N)
  begin
//    if (!Reset_N)             DataRdReady  <=  1'h0;
//    else 
    if (DataRdReadyClr)  DataRdReady  <=  1'h0;
    else if (DataRdEndReg)    DataRdReady  <=  1'h0;
    else if (DataRdEnd  )     DataRdReady  <=  1'h0;
    else if (DataRdEndFlag)   DataRdReady  <=  1'h0;
    else if (DataRdStart)     DataRdReady  <=  1'h1;
    else if (DataRdValid)     DataRdReady  <=  1'h1;
  end

  /////////////////////////////////////////////////////////

//22222222222222222222222222222222222222222222222222222




//3333333333333333333333333333333333333333333333333333333

  /////////////////////////////////////////////////////////
  wire [7:0]   RdByteNum =  AXI_BYTE_NUMBER ;
  reg  [31:0]  RdAddrCnt = 32'h0  ; //(O)[DdrRdCtrl]Ram Read Addrdss

  always @( posedge SysClk)
  begin
    if (DataRdStart)    RdAddrCnt <=  RdStartAddr;
    else  if (DataRdEn) RdAddrCnt <=  RdAddrCnt + {24'h0,RdByteNum};
  end

  /////////////////////////////////////////////////////////

  always @( posedge SysClk)   RamRdBusy <= DataRdReady | DataRdAddrAva;

  /////////////////////////////////////////////////////////
  reg   DataRdBusy = 1'h0;

  always @( posedge SysClk or negedge Reset_N)
  begin
  	if( !Reset_N ) 			DataRdBusy <=  1'h0;
    else if (DataRdEnd) DataRdBusy <=  1'h0;
    else if (DataRdEn)  DataRdBusy <=  1'h1;
  end

  /////////////////////////////////////////////////////////
  
  always @( posedge SysClk)  RamRdEnd  <=  DataRdEn & (~DataRdBusy) ;   //(O)[DdrRdCtrl]Ram Read End

  /////////////////////////////////////////////////////////
  
  always @( posedge SysClk)                 RamRdDAva <=  DataRdEn   ; //(O)[DdrRdCtrl]Ram Read Available
  always @( posedge SysClk)  if (DataRdEn)  RamRdData <=  DataRdData ; //(O)[DdrRdCtrl]Ram Read Data
  always @( posedge SysClk)  if (DataRdEn)  RamRdAddr <=  RdAddrCnt  ; //(O)[DdrRdCtrl]Ram Read Addrdss

//3333333333333333333333333333333333333333333333333333333

endmodule



